//******************************************
// Author: Jakub Zaroda
// Email: jakub.zaroda@outlook.com
//******************************************

module GiftPipeDecRoundFun(
    input wire inClk,
    input wire [127:0] inData,
    input wire [127:0] inKey,
    output wire [127:0] outData
);

wire [127:0] wireKey1;
wire [127:0] wireKey2;
wire [127:0] wireKey3;
wire [127:0] wireKey4;
wire [127:0] wireKey5;
wire [127:0] wireKey6;
wire [127:0] wireKey7;
wire [127:0] wireKey8;
wire [127:0] wireKey9;
wire [127:0] wireKey10;
wire [127:0] wireKey11;
wire [127:0] wireKey12;
wire [127:0] wireKey13;
wire [127:0] wireKey14;
wire [127:0] wireKey15;
wire [127:0] wireKey16;
wire [127:0] wireKey17;
wire [127:0] wireKey18;
wire [127:0] wireKey19;
wire [127:0] wireKey20;
wire [127:0] wireKey21;
wire [127:0] wireKey22;
wire [127:0] wireKey23;
wire [127:0] wireKey24;
wire [127:0] wireKey25;
wire [127:0] wireKey26;
wire [127:0] wireKey27;
wire [127:0] wireKey28;
wire [127:0] wireKey29;
wire [127:0] wireKey30;
wire [127:0] wireKey31;
wire [127:0] wireKey32;
wire [127:0] wireKey33;
wire [127:0] wireKey34;
wire [127:0] wireKey35;
wire [127:0] wireKey36;
wire [127:0] wireKey37;
wire [127:0] wireKey38;
wire [127:0] wireKey39;


wire [127:0] wireData1;
wire [127:0] wireData2;
wire [127:0] wireData3;
wire [127:0] wireData4;
wire [127:0] wireData5;
wire [127:0] wireData6;
wire [127:0] wireData7;
wire [127:0] wireData8;
wire [127:0] wireData9;
wire [127:0] wireData10;
wire [127:0] wireData11;
wire [127:0] wireData12;
wire [127:0] wireData13;
wire [127:0] wireData14;
wire [127:0] wireData15;
wire [127:0] wireData16;
wire [127:0] wireData17;
wire [127:0] wireData18;
wire [127:0] wireData19;
wire [127:0] wireData20;
wire [127:0] wireData21;
wire [127:0] wireData22;
wire [127:0] wireData23;
wire [127:0] wireData24;
wire [127:0] wireData25;
wire [127:0] wireData26;
wire [127:0] wireData27;
wire [127:0] wireData28;
wire [127:0] wireData29;
wire [127:0] wireData30;
wire [127:0] wireData31;
wire [127:0] wireData32;
wire [127:0] wireData33;
wire [127:0] wireData34;
wire [127:0] wireData35;
wire [127:0] wireData36;
wire [127:0] wireData37;
wire [127:0] wireData38;
wire [127:0] wireData39;


reg [127:0] regKey1 = 128'b0;
reg [127:0] regKey2 = 128'b0;
reg [127:0] regKey3 = 128'b0;
reg [127:0] regKey4 = 128'b0;
reg [127:0] regKey5 = 128'b0;
reg [127:0] regKey6 = 128'b0;
reg [127:0] regKey7 = 128'b0;
reg [127:0] regKey8 = 128'b0;
reg [127:0] regKey9 = 128'b0;
reg [127:0] regKey10 = 128'b0;
reg [127:0] regKey11 = 128'b0;
reg [127:0] regKey12 = 128'b0;
reg [127:0] regKey13 = 128'b0;
reg [127:0] regKey14 = 128'b0;
reg [127:0] regKey15 = 128'b0;
reg [127:0] regKey16 = 128'b0;
reg [127:0] regKey17 = 128'b0;
reg [127:0] regKey18 = 128'b0;
reg [127:0] regKey19 = 128'b0;
reg [127:0] regKey20 = 128'b0;
reg [127:0] regKey21 = 128'b0;
reg [127:0] regKey22 = 128'b0;
reg [127:0] regKey23 = 128'b0;
reg [127:0] regKey24 = 128'b0;
reg [127:0] regKey25 = 128'b0;
reg [127:0] regKey26 = 128'b0;
reg [127:0] regKey27 = 128'b0;
reg [127:0] regKey28 = 128'b0;
reg [127:0] regKey29 = 128'b0;
reg [127:0] regKey30 = 128'b0;
reg [127:0] regKey31 = 128'b0;
reg [127:0] regKey32 = 128'b0;
reg [127:0] regKey33 = 128'b0;
reg [127:0] regKey34 = 128'b0;
reg [127:0] regKey35 = 128'b0;
reg [127:0] regKey36 = 128'b0;
reg [127:0] regKey37 = 128'b0;
reg [127:0] regKey38 = 128'b0;
reg [127:0] regKey39 = 128'b0;
reg [127:0] regKey40 = 128'b0;

reg [5:0] regConstant1 = 6'h01;
reg [5:0] regConstant2 = 6'h03;
reg [5:0] regConstant3 = 6'h07;
reg [5:0] regConstant4 = 6'h0f;
reg [5:0] regConstant5 = 6'h1f;
reg [5:0] regConstant6 = 6'h3e;
reg [5:0] regConstant7 = 6'h3d;
reg [5:0] regConstant8 = 6'h3b;
reg [5:0] regConstant9 = 6'h37;
reg [5:0] regConstant10 = 6'h2f;
reg [5:0] regConstant11 = 6'h1e;
reg [5:0] regConstant12 = 6'h3c;
reg [5:0] regConstant13 = 6'h39;
reg [5:0] regConstant14 = 6'h33;
reg [5:0] regConstant15 = 6'h27;
reg [5:0] regConstant16 = 6'h0e;
reg [5:0] regConstant17 = 6'h1d;
reg [5:0] regConstant18 = 6'h3a;
reg [5:0] regConstant19 = 6'h35;
reg [5:0] regConstant20 = 6'h2b;
reg [5:0] regConstant21 = 6'h16;
reg [5:0] regConstant22 = 6'h2c;
reg [5:0] regConstant23 = 6'h18;
reg [5:0] regConstant24 = 6'h30;
reg [5:0] regConstant25 = 6'h21;
reg [5:0] regConstant26 = 6'h02;
reg [5:0] regConstant27 = 6'h05;
reg [5:0] regConstant28 = 6'h0b;
reg [5:0] regConstant29 = 6'h17;
reg [5:0] regConstant30 = 6'h2e;
reg [5:0] regConstant31 = 6'h1c;
reg [5:0] regConstant32 = 6'h38;
reg [5:0] regConstant33 = 6'h31;
reg [5:0] regConstant34 = 6'h23;
reg [5:0] regConstant35 = 6'h06;
reg [5:0] regConstant36 = 6'h0d;
reg [5:0] regConstant37 = 6'h1b;
reg [5:0] regConstant38 = 6'h36;
reg [5:0] regConstant39 = 6'h2d;
reg [5:0] regConstant40 = 6'h1a;


always @(posedge inClk) begin
    regKey1 <= inKey;
    regKey2 <= wireKey1;
    regKey3 <= wireKey2;
    regKey4 <= wireKey3;
    regKey5 <= wireKey4;
    regKey6 <= wireKey5;
    regKey7 <= wireKey6;
    regKey8 <= wireKey7;
    regKey9 <= wireKey8;
    regKey10 <= wireKey9;
    regKey11 <= wireKey10;
    regKey12 <= wireKey11;
    regKey13 <= wireKey12;
    regKey14 <= wireKey13;
    regKey15 <= wireKey14;
    regKey16 <= wireKey15;
    regKey17 <= wireKey16;
    regKey18 <= wireKey17;
    regKey19 <= wireKey18;
    regKey20 <= wireKey19;
    regKey21 <= wireKey20;
    regKey22 <= wireKey21;
    regKey23 <= wireKey22;
    regKey24 <= wireKey23;
    regKey25 <= wireKey24;
    regKey26 <= wireKey25;
    regKey27 <= wireKey26;
    regKey28 <= wireKey27;
    regKey29 <= wireKey28;
    regKey30 <= wireKey29;
    regKey31 <= wireKey30;
    regKey32 <= wireKey31;
    regKey33 <= wireKey32;
    regKey34 <= wireKey33;
    regKey35 <= wireKey34;
    regKey36 <= wireKey35;
    regKey37 <= wireKey36;
    regKey38 <= wireKey37;
    regKey39 <= wireKey38;
    regKey40 <= wireKey39;
end

GiftPipeInvKeyschFun instGiftPipeInvKeyschFun1 (.inData(regKey1), .outData(wireKey1));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun2 (.inData(regKey2), .outData(wireKey2));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun3 (.inData(regKey3), .outData(wireKey3));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun4 (.inData(regKey4), .outData(wireKey4));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun5 (.inData(regKey5), .outData(wireKey5));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun6 (.inData(regKey6), .outData(wireKey6));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun7 (.inData(regKey7), .outData(wireKey7));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun8 (.inData(regKey8), .outData(wireKey8));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun9 (.inData(regKey9), .outData(wireKey9));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun10 (.inData(regKey10), .outData(wireKey10));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun11 (.inData(regKey11), .outData(wireKey11));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun12 (.inData(regKey12), .outData(wireKey12));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun13 (.inData(regKey13), .outData(wireKey13));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun14 (.inData(regKey14), .outData(wireKey14));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun15 (.inData(regKey15), .outData(wireKey15));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun16 (.inData(regKey16), .outData(wireKey16));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun17 (.inData(regKey17), .outData(wireKey17));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun18 (.inData(regKey18), .outData(wireKey18));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun19 (.inData(regKey19), .outData(wireKey19));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun20 (.inData(regKey20), .outData(wireKey20));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun21 (.inData(regKey21), .outData(wireKey21));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun22 (.inData(regKey22), .outData(wireKey22));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun23 (.inData(regKey23), .outData(wireKey23));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun24 (.inData(regKey24), .outData(wireKey24));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun25 (.inData(regKey25), .outData(wireKey25));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun26 (.inData(regKey26), .outData(wireKey26));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun27 (.inData(regKey27), .outData(wireKey27));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun28 (.inData(regKey28), .outData(wireKey28));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun29 (.inData(regKey29), .outData(wireKey29));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun30 (.inData(regKey30), .outData(wireKey30));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun31 (.inData(regKey31), .outData(wireKey31));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun32 (.inData(regKey32), .outData(wireKey32));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun33 (.inData(regKey33), .outData(wireKey33));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun34 (.inData(regKey34), .outData(wireKey34));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun35 (.inData(regKey35), .outData(wireKey35));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun36 (.inData(regKey36), .outData(wireKey36));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun37 (.inData(regKey37), .outData(wireKey37));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun38 (.inData(regKey38), .outData(wireKey38));
GiftPipeInvKeyschFun instGiftPipeInvKeyschFun39 (.inData(regKey39), .outData(wireKey39));


reg [127:0] regData1 = 128'b0;
reg [127:0] regData2 = 128'b0;
reg [127:0] regData3 = 128'b0;
reg [127:0] regData4 = 128'b0;
reg [127:0] regData5 = 128'b0;
reg [127:0] regData6 = 128'b0;
reg [127:0] regData7 = 128'b0;
reg [127:0] regData8 = 128'b0;
reg [127:0] regData9 = 128'b0;
reg [127:0] regData10 = 128'b0;
reg [127:0] regData11 = 128'b0;
reg [127:0] regData12 = 128'b0;
reg [127:0] regData13 = 128'b0;
reg [127:0] regData14 = 128'b0;
reg [127:0] regData15 = 128'b0;
reg [127:0] regData16 = 128'b0;
reg [127:0] regData17 = 128'b0;
reg [127:0] regData18 = 128'b0;
reg [127:0] regData19 = 128'b0;
reg [127:0] regData20 = 128'b0;
reg [127:0] regData21 = 128'b0;
reg [127:0] regData22 = 128'b0;
reg [127:0] regData23 = 128'b0;
reg [127:0] regData24 = 128'b0;
reg [127:0] regData25 = 128'b0;
reg [127:0] regData26 = 128'b0;
reg [127:0] regData27 = 128'b0;
reg [127:0] regData28 = 128'b0;
reg [127:0] regData29 = 128'b0;
reg [127:0] regData30 = 128'b0;
reg [127:0] regData31 = 128'b0;
reg [127:0] regData32 = 128'b0;
reg [127:0] regData33 = 128'b0;
reg [127:0] regData34 = 128'b0;
reg [127:0] regData35 = 128'b0;
reg [127:0] regData36 = 128'b0;
reg [127:0] regData37 = 128'b0;
reg [127:0] regData38 = 128'b0;
reg [127:0] regData39 = 128'b0;
reg [127:0] regData40 = 128'b0;

always @(posedge inClk ) begin
    regData1 <= inData;
    regData2 <= wireData1;
    regData3 <= wireData2;
    regData4 <= wireData3;
    regData5 <= wireData4;
    regData6 <= wireData5;
    regData7 <= wireData6;
    regData8 <= wireData7;
    regData9 <= wireData8;
    regData10 <= wireData9;
    regData11 <= wireData10;
    regData12 <= wireData11;
    regData13 <= wireData12;
    regData14 <= wireData13;
    regData15 <= wireData14;
    regData16 <= wireData15;
    regData17 <= wireData16;
    regData18 <= wireData17;
    regData19 <= wireData18;
    regData20 <= wireData19;
    regData21 <= wireData20;
    regData22 <= wireData21;
    regData23 <= wireData22;
    regData24 <= wireData23;
    regData25 <= wireData24;
    regData26 <= wireData25;
    regData27 <= wireData26;
    regData28 <= wireData27;
    regData29 <= wireData28;
    regData30 <= wireData29;
    regData31 <= wireData30;
    regData32 <= wireData31;
    regData33 <= wireData32;
    regData34 <= wireData33;
    regData35 <= wireData34;
    regData36 <= wireData35;
    regData37 <= wireData36;
    regData38 <= wireData37;
    regData39 <= wireData38;
    regData40 <= wireData39;
end




GiftFullInvRoundFun instGiftFullInvRoundFun0 (.inData(regData1), .inKey(regKey1), .inConstant(regConstant40), .outData(wireData1));
GiftFullInvRoundFun instGiftFullInvRoundFun1 (.inData(regData2), .inKey(regKey2), .inConstant(regConstant39), .outData(wireData2));
GiftFullInvRoundFun instGiftFullInvRoundFun2 (.inData(regData3), .inKey(regKey3), .inConstant(regConstant38), .outData(wireData3));
GiftFullInvRoundFun instGiftFullInvRoundFun3 (.inData(regData4), .inKey(regKey4), .inConstant(regConstant37), .outData(wireData4));
GiftFullInvRoundFun instGiftFullInvRoundFun4 (.inData(regData5), .inKey(regKey5), .inConstant(regConstant36), .outData(wireData5));
GiftFullInvRoundFun instGiftFullInvRoundFun5 (.inData(regData6), .inKey(regKey6), .inConstant(regConstant35), .outData(wireData6));
GiftFullInvRoundFun instGiftFullInvRoundFun6 (.inData(regData7), .inKey(regKey7), .inConstant(regConstant34), .outData(wireData7));
GiftFullInvRoundFun instGiftFullInvRoundFun7 (.inData(regData8), .inKey(regKey8), .inConstant(regConstant33), .outData(wireData8));
GiftFullInvRoundFun instGiftFullInvRoundFun8 (.inData(regData9), .inKey(regKey9), .inConstant(regConstant32), .outData(wireData9));
GiftFullInvRoundFun instGiftFullInvRoundFun9 (.inData(regData10), .inKey(regKey10), .inConstant(regConstant31), .outData(wireData10));
GiftFullInvRoundFun instGiftFullInvRoundFun10 (.inData(regData11), .inKey(regKey11), .inConstant(regConstant30), .outData(wireData11));
GiftFullInvRoundFun instGiftFullInvRoundFun11 (.inData(regData12), .inKey(regKey12), .inConstant(regConstant29), .outData(wireData12));
GiftFullInvRoundFun instGiftFullInvRoundFun12 (.inData(regData13), .inKey(regKey13), .inConstant(regConstant28), .outData(wireData13));
GiftFullInvRoundFun instGiftFullInvRoundFun13 (.inData(regData14), .inKey(regKey14), .inConstant(regConstant27), .outData(wireData14));
GiftFullInvRoundFun instGiftFullInvRoundFun14 (.inData(regData15), .inKey(regKey15), .inConstant(regConstant26), .outData(wireData15));
GiftFullInvRoundFun instGiftFullInvRoundFun15 (.inData(regData16), .inKey(regKey16), .inConstant(regConstant25), .outData(wireData16));
GiftFullInvRoundFun instGiftFullInvRoundFun16 (.inData(regData17), .inKey(regKey17), .inConstant(regConstant24), .outData(wireData17));
GiftFullInvRoundFun instGiftFullInvRoundFun17 (.inData(regData18), .inKey(regKey18), .inConstant(regConstant23), .outData(wireData18));
GiftFullInvRoundFun instGiftFullInvRoundFun18 (.inData(regData19), .inKey(regKey19), .inConstant(regConstant22), .outData(wireData19));
GiftFullInvRoundFun instGiftFullInvRoundFun19 (.inData(regData20), .inKey(regKey20), .inConstant(regConstant21), .outData(wireData20));
GiftFullInvRoundFun instGiftFullInvRoundFun20 (.inData(regData21), .inKey(regKey21), .inConstant(regConstant20), .outData(wireData21));
GiftFullInvRoundFun instGiftFullInvRoundFun21 (.inData(regData22), .inKey(regKey22), .inConstant(regConstant19), .outData(wireData22));
GiftFullInvRoundFun instGiftFullInvRoundFun22 (.inData(regData23), .inKey(regKey23), .inConstant(regConstant18), .outData(wireData23));
GiftFullInvRoundFun instGiftFullInvRoundFun23 (.inData(regData24), .inKey(regKey24), .inConstant(regConstant17), .outData(wireData24));
GiftFullInvRoundFun instGiftFullInvRoundFun24 (.inData(regData25), .inKey(regKey25), .inConstant(regConstant16), .outData(wireData25));
GiftFullInvRoundFun instGiftFullInvRoundFun25 (.inData(regData26), .inKey(regKey26), .inConstant(regConstant15), .outData(wireData26));
GiftFullInvRoundFun instGiftFullInvRoundFun26 (.inData(regData27), .inKey(regKey27), .inConstant(regConstant14), .outData(wireData27));
GiftFullInvRoundFun instGiftFullInvRoundFun27 (.inData(regData28), .inKey(regKey28), .inConstant(regConstant13), .outData(wireData28));
GiftFullInvRoundFun instGiftFullInvRoundFun28 (.inData(regData29), .inKey(regKey29), .inConstant(regConstant12), .outData(wireData29));
GiftFullInvRoundFun instGiftFullInvRoundFun29 (.inData(regData30), .inKey(regKey30), .inConstant(regConstant11), .outData(wireData30));
GiftFullInvRoundFun instGiftFullInvRoundFun30 (.inData(regData31), .inKey(regKey31), .inConstant(regConstant10), .outData(wireData31));
GiftFullInvRoundFun instGiftFullInvRoundFun31 (.inData(regData32), .inKey(regKey32), .inConstant(regConstant9), .outData(wireData32));
GiftFullInvRoundFun instGiftFullInvRoundFun32 (.inData(regData33), .inKey(regKey33), .inConstant(regConstant8), .outData(wireData33));
GiftFullInvRoundFun instGiftFullInvRoundFun33 (.inData(regData34), .inKey(regKey34), .inConstant(regConstant7), .outData(wireData34));
GiftFullInvRoundFun instGiftFullInvRoundFun34 (.inData(regData35), .inKey(regKey35), .inConstant(regConstant6), .outData(wireData35));
GiftFullInvRoundFun instGiftFullInvRoundFun35 (.inData(regData36), .inKey(regKey36), .inConstant(regConstant5), .outData(wireData36));
GiftFullInvRoundFun instGiftFullInvRoundFun36 (.inData(regData37), .inKey(regKey37), .inConstant(regConstant4), .outData(wireData37));
GiftFullInvRoundFun instGiftFullInvRoundFun37 (.inData(regData38), .inKey(regKey38), .inConstant(regConstant3), .outData(wireData38));
GiftFullInvRoundFun instGiftFullInvRoundFun38 (.inData(regData39), .inKey(regKey39), .inConstant(regConstant2), .outData(wireData39));
GiftFullInvRoundFun instGiftFullInvRoundFun39 (.inData(regData40), .inKey(regKey40), .inConstant(regConstant1), .outData(outData));



endmodule