//******************************************
// Author: Jakub Zaroda
// Email: jakub.zaroda@outlook.com
//******************************************

module GiftFullRoundFun(
    input wire [127:0] inData,
    input wire [127:0] inKey,
    input wire [5:0]   inConstant,
    output wire [127:0] outData
);

wire [127:0] wireKey1;
wire [127:0] wireKey2;
wire [127:0] wireKey3;
wire [127:0] wireKey4;
wire [127:0] wireKey5;
wire [127:0] wireKey6;
wire [127:0] wireKey7;
wire [127:0] wireKey8;
wire [127:0] wireKey9;
wire [127:0] wireKey10;
wire [127:0] wireKey11;
wire [127:0] wireKey12;
wire [127:0] wireKey13;
wire [127:0] wireKey14;
wire [127:0] wireKey15;
wire [127:0] wireKey16;
wire [127:0] wireKey17;
wire [127:0] wireKey18;
wire [127:0] wireKey19;
wire [127:0] wireKey20;
wire [127:0] wireKey21;
wire [127:0] wireKey22;
wire [127:0] wireKey23;
wire [127:0] wireKey24;
wire [127:0] wireKey25;
wire [127:0] wireKey26;
wire [127:0] wireKey27;
wire [127:0] wireKey28;
wire [127:0] wireKey29;
wire [127:0] wireKey30;
wire [127:0] wireKey31;
wire [127:0] wireKey32;
wire [127:0] wireKey33;
wire [127:0] wireKey34;
wire [127:0] wireKey35;
wire [127:0] wireKey36;
wire [127:0] wireKey37;
wire [127:0] wireKey38;
wire [127:0] wireKey39;

wire [5:0] wireConstant1;
wire [5:0] wireConstant2;
wire [5:0] wireConstant3;
wire [5:0] wireConstant4;
wire [5:0] wireConstant5;
wire [5:0] wireConstant6;
wire [5:0] wireConstant7;
wire [5:0] wireConstant8;
wire [5:0] wireConstant9;
wire [5:0] wireConstant10;
wire [5:0] wireConstant11;
wire [5:0] wireConstant12;
wire [5:0] wireConstant13;
wire [5:0] wireConstant14;
wire [5:0] wireConstant15;
wire [5:0] wireConstant16;
wire [5:0] wireConstant17;
wire [5:0] wireConstant18;
wire [5:0] wireConstant19;
wire [5:0] wireConstant20;
wire [5:0] wireConstant21;
wire [5:0] wireConstant22;
wire [5:0] wireConstant23;
wire [5:0] wireConstant24;
wire [5:0] wireConstant25;
wire [5:0] wireConstant26;
wire [5:0] wireConstant27;
wire [5:0] wireConstant28;
wire [5:0] wireConstant29;
wire [5:0] wireConstant30;
wire [5:0] wireConstant31;
wire [5:0] wireConstant32;
wire [5:0] wireConstant33;
wire [5:0] wireConstant34;
wire [5:0] wireConstant35;
wire [5:0] wireConstant36;
wire [5:0] wireConstant37;
wire [5:0] wireConstant38;
wire [5:0] wireConstant39;

wire [127:0] wireData1;
wire [127:0] wireData2;
wire [127:0] wireData3;
wire [127:0] wireData4;
wire [127:0] wireData5;
wire [127:0] wireData6;
wire [127:0] wireData7;
wire [127:0] wireData8;
wire [127:0] wireData9;
wire [127:0] wireData10;
wire [127:0] wireData11;
wire [127:0] wireData12;
wire [127:0] wireData13;
wire [127:0] wireData14;
wire [127:0] wireData15;
wire [127:0] wireData16;
wire [127:0] wireData17;
wire [127:0] wireData18;
wire [127:0] wireData19;
wire [127:0] wireData20;
wire [127:0] wireData21;
wire [127:0] wireData22;
wire [127:0] wireData23;
wire [127:0] wireData24;
wire [127:0] wireData25;
wire [127:0] wireData26;
wire [127:0] wireData27;
wire [127:0] wireData28;
wire [127:0] wireData29;
wire [127:0] wireData30;
wire [127:0] wireData31;
wire [127:0] wireData32;
wire [127:0] wireData33;
wire [127:0] wireData34;
wire [127:0] wireData35;
wire [127:0] wireData36;
wire [127:0] wireData37;
wire [127:0] wireData38;
wire [127:0] wireData39;


GiftKeyschFun instGiftKeyschFun1 (.inData(inKey), .outData(wireKey1));
GiftKeyschFun instGiftKeyschFun2 (.inData(wireKey1), .outData(wireKey2));
GiftKeyschFun instGiftKeyschFun3 (.inData(wireKey2), .outData(wireKey3));
GiftKeyschFun instGiftKeyschFun4 (.inData(wireKey3), .outData(wireKey4));
GiftKeyschFun instGiftKeyschFun5 (.inData(wireKey4), .outData(wireKey5));
GiftKeyschFun instGiftKeyschFun6 (.inData(wireKey5), .outData(wireKey6));
GiftKeyschFun instGiftKeyschFun7 (.inData(wireKey6), .outData(wireKey7));
GiftKeyschFun instGiftKeyschFun8 (.inData(wireKey7), .outData(wireKey8));
GiftKeyschFun instGiftKeyschFun9 (.inData(wireKey8), .outData(wireKey9));
GiftKeyschFun instGiftKeyschFun10 (.inData(wireKey9), .outData(wireKey10));
GiftKeyschFun instGiftKeyschFun11 (.inData(wireKey10), .outData(wireKey11));
GiftKeyschFun instGiftKeyschFun12 (.inData(wireKey11), .outData(wireKey12));
GiftKeyschFun instGiftKeyschFun13 (.inData(wireKey12), .outData(wireKey13));
GiftKeyschFun instGiftKeyschFun14 (.inData(wireKey13), .outData(wireKey14));
GiftKeyschFun instGiftKeyschFun15 (.inData(wireKey14), .outData(wireKey15));
GiftKeyschFun instGiftKeyschFun16 (.inData(wireKey15), .outData(wireKey16));
GiftKeyschFun instGiftKeyschFun17 (.inData(wireKey16), .outData(wireKey17));
GiftKeyschFun instGiftKeyschFun18 (.inData(wireKey17), .outData(wireKey18));
GiftKeyschFun instGiftKeyschFun19 (.inData(wireKey18), .outData(wireKey19));
GiftKeyschFun instGiftKeyschFun20 (.inData(wireKey19), .outData(wireKey20));
GiftKeyschFun instGiftKeyschFun21 (.inData(wireKey20), .outData(wireKey21));
GiftKeyschFun instGiftKeyschFun22 (.inData(wireKey21), .outData(wireKey22));
GiftKeyschFun instGiftKeyschFun23 (.inData(wireKey22), .outData(wireKey23));
GiftKeyschFun instGiftKeyschFun24 (.inData(wireKey23), .outData(wireKey24));
GiftKeyschFun instGiftKeyschFun25 (.inData(wireKey24), .outData(wireKey25));
GiftKeyschFun instGiftKeyschFun26 (.inData(wireKey25), .outData(wireKey26));
GiftKeyschFun instGiftKeyschFun27 (.inData(wireKey26), .outData(wireKey27));
GiftKeyschFun instGiftKeyschFun28 (.inData(wireKey27), .outData(wireKey28));
GiftKeyschFun instGiftKeyschFun29 (.inData(wireKey28), .outData(wireKey29));
GiftKeyschFun instGiftKeyschFun30 (.inData(wireKey29), .outData(wireKey30));
GiftKeyschFun instGiftKeyschFun31 (.inData(wireKey30), .outData(wireKey31));
GiftKeyschFun instGiftKeyschFun32 (.inData(wireKey31), .outData(wireKey32));
GiftKeyschFun instGiftKeyschFun33 (.inData(wireKey32), .outData(wireKey33));
GiftKeyschFun instGiftKeyschFun34 (.inData(wireKey33), .outData(wireKey34));
GiftKeyschFun instGiftKeyschFun35 (.inData(wireKey34), .outData(wireKey35));
GiftKeyschFun instGiftKeyschFun36 (.inData(wireKey35), .outData(wireKey36));
GiftKeyschFun instGiftKeyschFun37 (.inData(wireKey36), .outData(wireKey37));
GiftKeyschFun instGiftKeyschFun38 (.inData(wireKey37), .outData(wireKey38));
GiftKeyschFun instGiftKeyschFun39 (.inData(wireKey38), .outData(wireKey39));

GiftConstFun instGiftConstFun1 (.inData(inConstant), .outData(wireConstant1));
GiftConstFun instGiftConstFun2 (.inData(wireConstant1), .outData(wireConstant2));
GiftConstFun instGiftConstFun3 (.inData(wireConstant2), .outData(wireConstant3));
GiftConstFun instGiftConstFun4 (.inData(wireConstant3), .outData(wireConstant4));
GiftConstFun instGiftConstFun5 (.inData(wireConstant4), .outData(wireConstant5));
GiftConstFun instGiftConstFun6 (.inData(wireConstant5), .outData(wireConstant6));
GiftConstFun instGiftConstFun7 (.inData(wireConstant6), .outData(wireConstant7));
GiftConstFun instGiftConstFun8 (.inData(wireConstant7), .outData(wireConstant8));
GiftConstFun instGiftConstFun9 (.inData(wireConstant8), .outData(wireConstant9));
GiftConstFun instGiftConstFun10 (.inData(wireConstant9), .outData(wireConstant10));
GiftConstFun instGiftConstFun11 (.inData(wireConstant10), .outData(wireConstant11));
GiftConstFun instGiftConstFun12 (.inData(wireConstant11), .outData(wireConstant12));
GiftConstFun instGiftConstFun13 (.inData(wireConstant12), .outData(wireConstant13));
GiftConstFun instGiftConstFun14 (.inData(wireConstant13), .outData(wireConstant14));
GiftConstFun instGiftConstFun15 (.inData(wireConstant14), .outData(wireConstant15));
GiftConstFun instGiftConstFun16 (.inData(wireConstant15), .outData(wireConstant16));
GiftConstFun instGiftConstFun17 (.inData(wireConstant16), .outData(wireConstant17));
GiftConstFun instGiftConstFun18 (.inData(wireConstant17), .outData(wireConstant18));
GiftConstFun instGiftConstFun19 (.inData(wireConstant18), .outData(wireConstant19));
GiftConstFun instGiftConstFun20 (.inData(wireConstant19), .outData(wireConstant20));
GiftConstFun instGiftConstFun21 (.inData(wireConstant20), .outData(wireConstant21));
GiftConstFun instGiftConstFun22 (.inData(wireConstant21), .outData(wireConstant22));
GiftConstFun instGiftConstFun23 (.inData(wireConstant22), .outData(wireConstant23));
GiftConstFun instGiftConstFun24 (.inData(wireConstant23), .outData(wireConstant24));
GiftConstFun instGiftConstFun25 (.inData(wireConstant24), .outData(wireConstant25));
GiftConstFun instGiftConstFun26 (.inData(wireConstant25), .outData(wireConstant26));
GiftConstFun instGiftConstFun27 (.inData(wireConstant26), .outData(wireConstant27));
GiftConstFun instGiftConstFun28 (.inData(wireConstant27), .outData(wireConstant28));
GiftConstFun instGiftConstFun29 (.inData(wireConstant28), .outData(wireConstant29));
GiftConstFun instGiftConstFun30 (.inData(wireConstant29), .outData(wireConstant30));
GiftConstFun instGiftConstFun31 (.inData(wireConstant30), .outData(wireConstant31));
GiftConstFun instGiftConstFun32 (.inData(wireConstant31), .outData(wireConstant32));
GiftConstFun instGiftConstFun33 (.inData(wireConstant32), .outData(wireConstant33));
GiftConstFun instGiftConstFun34 (.inData(wireConstant33), .outData(wireConstant34));
GiftConstFun instGiftConstFun35 (.inData(wireConstant34), .outData(wireConstant35));
GiftConstFun instGiftConstFun36 (.inData(wireConstant35), .outData(wireConstant36));
GiftConstFun instGiftConstFun37 (.inData(wireConstant36), .outData(wireConstant37));
GiftConstFun instGiftConstFun38 (.inData(wireConstant37), .outData(wireConstant38));
GiftConstFun instGiftConstFun39 (.inData(wireConstant38), .outData(wireConstant39));



GiftRoundFun instGiftRoundFun0 (.inData(inData), .inKey(inKey), .inConstant(inConstant), .outData(wireData1));
GiftRoundFun instGiftRoundFun1 (.inData(wireData1), .inKey(wireKey1), .inConstant(wireConstant1), .outData(wireData2));
GiftRoundFun instGiftRoundFun2 (.inData(wireData2), .inKey(wireKey2), .inConstant(wireConstant2), .outData(wireData3));
GiftRoundFun instGiftRoundFun3 (.inData(wireData3), .inKey(wireKey3), .inConstant(wireConstant3), .outData(wireData4));
GiftRoundFun instGiftRoundFun4 (.inData(wireData4), .inKey(wireKey4), .inConstant(wireConstant4), .outData(wireData5));
GiftRoundFun instGiftRoundFun5 (.inData(wireData5), .inKey(wireKey5), .inConstant(wireConstant5), .outData(wireData6));
GiftRoundFun instGiftRoundFun6 (.inData(wireData6), .inKey(wireKey6), .inConstant(wireConstant6), .outData(wireData7));
GiftRoundFun instGiftRoundFun7 (.inData(wireData7), .inKey(wireKey7), .inConstant(wireConstant7), .outData(wireData8));
GiftRoundFun instGiftRoundFun8 (.inData(wireData8), .inKey(wireKey8), .inConstant(wireConstant8), .outData(wireData9));
GiftRoundFun instGiftRoundFun9 (.inData(wireData9), .inKey(wireKey9), .inConstant(wireConstant9), .outData(wireData10));
GiftRoundFun instGiftRoundFun10 (.inData(wireData10), .inKey(wireKey10), .inConstant(wireConstant10), .outData(wireData11));
GiftRoundFun instGiftRoundFun11 (.inData(wireData11), .inKey(wireKey11), .inConstant(wireConstant11), .outData(wireData12));
GiftRoundFun instGiftRoundFun12 (.inData(wireData12), .inKey(wireKey12), .inConstant(wireConstant12), .outData(wireData13));
GiftRoundFun instGiftRoundFun13 (.inData(wireData13), .inKey(wireKey13), .inConstant(wireConstant13), .outData(wireData14));
GiftRoundFun instGiftRoundFun14 (.inData(wireData14), .inKey(wireKey14), .inConstant(wireConstant14), .outData(wireData15));
GiftRoundFun instGiftRoundFun15 (.inData(wireData15), .inKey(wireKey15), .inConstant(wireConstant15), .outData(wireData16));
GiftRoundFun instGiftRoundFun16 (.inData(wireData16), .inKey(wireKey16), .inConstant(wireConstant16), .outData(wireData17));
GiftRoundFun instGiftRoundFun17 (.inData(wireData17), .inKey(wireKey17), .inConstant(wireConstant17), .outData(wireData18));
GiftRoundFun instGiftRoundFun18 (.inData(wireData18), .inKey(wireKey18), .inConstant(wireConstant18), .outData(wireData19));
GiftRoundFun instGiftRoundFun19 (.inData(wireData19), .inKey(wireKey19), .inConstant(wireConstant19), .outData(wireData20));
GiftRoundFun instGiftRoundFun20 (.inData(wireData20), .inKey(wireKey20), .inConstant(wireConstant20), .outData(wireData21));
GiftRoundFun instGiftRoundFun21 (.inData(wireData21), .inKey(wireKey21), .inConstant(wireConstant21), .outData(wireData22));
GiftRoundFun instGiftRoundFun22 (.inData(wireData22), .inKey(wireKey22), .inConstant(wireConstant22), .outData(wireData23));
GiftRoundFun instGiftRoundFun23 (.inData(wireData23), .inKey(wireKey23), .inConstant(wireConstant23), .outData(wireData24));
GiftRoundFun instGiftRoundFun24 (.inData(wireData24), .inKey(wireKey24), .inConstant(wireConstant24), .outData(wireData25));
GiftRoundFun instGiftRoundFun25 (.inData(wireData25), .inKey(wireKey25), .inConstant(wireConstant25), .outData(wireData26));
GiftRoundFun instGiftRoundFun26 (.inData(wireData26), .inKey(wireKey26), .inConstant(wireConstant26), .outData(wireData27));
GiftRoundFun instGiftRoundFun27 (.inData(wireData27), .inKey(wireKey27), .inConstant(wireConstant27), .outData(wireData28));
GiftRoundFun instGiftRoundFun28 (.inData(wireData28), .inKey(wireKey28), .inConstant(wireConstant28), .outData(wireData29));
GiftRoundFun instGiftRoundFun29 (.inData(wireData29), .inKey(wireKey29), .inConstant(wireConstant29), .outData(wireData30));
GiftRoundFun instGiftRoundFun30 (.inData(wireData30), .inKey(wireKey30), .inConstant(wireConstant30), .outData(wireData31));
GiftRoundFun instGiftRoundFun31 (.inData(wireData31), .inKey(wireKey31), .inConstant(wireConstant31), .outData(wireData32));
GiftRoundFun instGiftRoundFun32 (.inData(wireData32), .inKey(wireKey32), .inConstant(wireConstant32), .outData(wireData33));
GiftRoundFun instGiftRoundFun33 (.inData(wireData33), .inKey(wireKey33), .inConstant(wireConstant33), .outData(wireData34));
GiftRoundFun instGiftRoundFun34 (.inData(wireData34), .inKey(wireKey34), .inConstant(wireConstant34), .outData(wireData35));
GiftRoundFun instGiftRoundFun35 (.inData(wireData35), .inKey(wireKey35), .inConstant(wireConstant35), .outData(wireData36));
GiftRoundFun instGiftRoundFun36 (.inData(wireData36), .inKey(wireKey36), .inConstant(wireConstant36), .outData(wireData37));
GiftRoundFun instGiftRoundFun37 (.inData(wireData37), .inKey(wireKey37), .inConstant(wireConstant37), .outData(wireData38));
GiftRoundFun instGiftRoundFun38 (.inData(wireData38), .inKey(wireKey38), .inConstant(wireConstant38), .outData(wireData39));
GiftRoundFun instGiftRoundFun39 (.inData(wireData39), .inKey(wireKey39), .inConstant(wireConstant39), .outData(outData));



endmodule