//******************************************
// Author: Jakub Zaroda
// Email: jakub.zaroda@outlook.com
//******************************************

module GiftPermutationFun (
    input wire [127:0] inData,
    output wire [127:0] outData
);

assign outData[0] = inData[0];
assign outData[33] = inData[1];
assign outData[66] = inData[2];
assign outData[99] = inData[3];
assign outData[96] = inData[4];
assign outData[1] = inData[5];
assign outData[34] = inData[6];
assign outData[67] = inData[7];
assign outData[64] = inData[8];
assign outData[97] = inData[9];
assign outData[2] = inData[10];
assign outData[35] = inData[11];
assign outData[32] = inData[12];
assign outData[65] = inData[13];
assign outData[98] = inData[14];
assign outData[3] = inData[15];
assign outData[4] = inData[16];
assign outData[37] = inData[17];
assign outData[70] = inData[18];
assign outData[103] = inData[19];
assign outData[100] = inData[20];
assign outData[5] = inData[21];
assign outData[38] = inData[22];
assign outData[71] = inData[23];
assign outData[68] = inData[24];
assign outData[101] = inData[25];
assign outData[6] = inData[26];
assign outData[39] = inData[27];
assign outData[36] = inData[28];
assign outData[69] = inData[29];
assign outData[102] = inData[30];
assign outData[7] = inData[31];
assign outData[8] = inData[32];
assign outData[41] = inData[33];
assign outData[74] = inData[34];
assign outData[107] = inData[35];
assign outData[104] = inData[36];
assign outData[9] = inData[37];
assign outData[42] = inData[38];
assign outData[75] = inData[39];
assign outData[72] = inData[40];
assign outData[105] = inData[41];
assign outData[10] = inData[42];
assign outData[43] = inData[43];
assign outData[40] = inData[44];
assign outData[73] = inData[45];
assign outData[106] = inData[46];
assign outData[11] = inData[47];
assign outData[12] = inData[48];
assign outData[45] = inData[49];
assign outData[78] = inData[50];
assign outData[111] = inData[51];
assign outData[108] = inData[52];
assign outData[13] = inData[53];
assign outData[46] = inData[54];
assign outData[79] = inData[55];
assign outData[76] = inData[56];
assign outData[109] = inData[57];
assign outData[14] = inData[58];
assign outData[47] = inData[59];
assign outData[44] = inData[60];
assign outData[77] = inData[61];
assign outData[110] = inData[62];
assign outData[15] = inData[63];
assign outData[16] = inData[64];
assign outData[49] = inData[65];
assign outData[82] = inData[66];
assign outData[115] = inData[67];
assign outData[112] = inData[68];
assign outData[17] = inData[69];
assign outData[50] = inData[70];
assign outData[83] = inData[71];
assign outData[80] = inData[72];
assign outData[113] = inData[73];
assign outData[18] = inData[74];
assign outData[51] = inData[75];
assign outData[48] = inData[76];
assign outData[81] = inData[77];
assign outData[114] = inData[78];
assign outData[19] = inData[79];
assign outData[20] = inData[80];
assign outData[53] = inData[81];
assign outData[86] = inData[82];
assign outData[119] = inData[83];
assign outData[116] = inData[84];
assign outData[21] = inData[85];
assign outData[54] = inData[86];
assign outData[87] = inData[87];
assign outData[84] = inData[88];
assign outData[117] = inData[89];
assign outData[22] = inData[90];
assign outData[55] = inData[91];
assign outData[52] = inData[92];
assign outData[85] = inData[93];
assign outData[118] = inData[94];
assign outData[23] = inData[95];
assign outData[24] = inData[96];
assign outData[57] = inData[97];
assign outData[90] = inData[98];
assign outData[123] = inData[99];
assign outData[120] = inData[100];
assign outData[25] = inData[101];
assign outData[58] = inData[102];
assign outData[91] = inData[103];
assign outData[88] = inData[104];
assign outData[121] = inData[105];
assign outData[26] = inData[106];
assign outData[59] = inData[107];
assign outData[56] = inData[108];
assign outData[89] = inData[109];
assign outData[122] = inData[110];
assign outData[27] = inData[111];
assign outData[28] = inData[112];
assign outData[61] = inData[113];
assign outData[94] = inData[114];
assign outData[127] = inData[115];
assign outData[124] = inData[116];
assign outData[29] = inData[117];
assign outData[62] = inData[118];
assign outData[95] = inData[119];
assign outData[92] = inData[120];
assign outData[125] = inData[121];
assign outData[30] = inData[122];
assign outData[63] = inData[123];
assign outData[60] = inData[124];
assign outData[93] = inData[125];
assign outData[126] = inData[126];
assign outData[31] = inData[127];

endmodule